library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity full_adder is
    Port ( a,b : in std_logic;
           c : out std_logic);
end full_adder;

architecture Behavioral of full_adder is

begin


end Behavioral;
